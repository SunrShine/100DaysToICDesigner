module ringCounter(
    port_list
);
    
endmodule