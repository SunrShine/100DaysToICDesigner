module tester(model1_bfm bfm);


endmodule