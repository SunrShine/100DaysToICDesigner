module Sync_fifo #(parameter WIDTH = 8) (
    input wire clk,
    input wire rst_n,

);
    
endmodule                                                                                                                                                                                                                                                                                                                                                                    