module tb_fdiv8_7;


endmodule //tb_fdiv8_7