module Decoder_4_16 (
    ports
);
    
endmodule