module top();
    
    
endmodule