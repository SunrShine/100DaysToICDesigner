module tb_ahb_master_port;



endmodule