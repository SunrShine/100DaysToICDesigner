module DLatch (
    input wire R,  //复位
    input wire S,   //置位
    input wire C,  //使能
    output reg Q,
    output reg Q_n
);
    


endmodule

