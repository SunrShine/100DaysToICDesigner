module lookaheadCarryAdder #(
    parameters width = 4
) (
    ports
);
    //超前进位加法器的思想是并行计算进位, 
    //通过公式直接导出最终结果与每个输入的关系,
    //是一种用面积换性能的方法



endmodule



//子模块，计算进位
