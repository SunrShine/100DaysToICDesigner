
package xpk;
    int x;
    class x1;
        
    endclass
endpackage

package A;
    import xpk::x1;
    int b;
    class A1 extends x1;
        
    endclass

endpackage

package B;
    
    
endpackage