module divthree(
    input wire clk,
    input wire rst_n,
    
);
    
endmodule