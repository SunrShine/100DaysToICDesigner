module tb_autosale;
    
endmodule